class asyn_fifo_base_read_sequence extends uvm_sequence #(asyn_fifo_read_sequence_item);
	`uvm_object_utils(asyn_fifo_base_read_sequence)

	function new(string name = "asyn_fifo_base_read_sequence");
		super.new(name);
	endfunction

	virtual task body();
		req = asyn_fifo_read_sequence_item::type_id::create("req");
		wait_for_grant();
		req.randomize();
		send_request(req);
		wait_for_item_done();
	endtask
endclass
//-------------------------------------------------------------------------------------------------------------------
// Read Reset Sequence
//-------------------------------------------------------------------------------------------------------------------
class read_reset_sequence extends uvm_sequence #(asyn_fifo_read_sequence_item); 
		`uvm_object_utils(read_reset_sequence)

		function new(string name = "read_reset_sequence");
			super.new(name);
		endfunction

		virtual task body();
			`uvm_do_with(req,{req.rrst_n == 'b0;});
		endtask
endclass
