`include "uvm_macros.svh"
package asyn_fifo_pkg;
	`include "asyn_fifo_write_sequence_item.sv"
	`include "asyn_fifo_read_sequence_item.sv"

	`include "asyn_fifo_write_sequencer.sv"
	`include "asyn_fifo_read_sequencer.sv"

	`include "asyn_fifo_write_sequence.sv"
	`include "asyn_fifo_read_sequence.sv"

	`include "asyn_fifo_virtual_sequencer.sv"
	`include "asyn_fifo_virtual_sequence.sv"
	`include "asyn_fifo_write_driver.sv"
	`include "asyn_fifo_read_driver.sv"
	`include "asyn_fifo_write_monitor.sv"
	`include "asyn_fifo_read_monitor.sv"
	`include "asyn_fifo_write_agent.sv"
	`include "asyn_fifo_read_agent.sv"
	`include "asyn_fifo_scoreboard.sv"
	`include "asyn_fifo_subscriber.sv"
	`include "asyn_fifo_env.sv"
	`include "asyn_fifo_test.sv"
endpackage
