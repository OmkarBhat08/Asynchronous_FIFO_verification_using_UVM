`define DSIZE 8
`define A_SIZE 4
